module mixer(
	input wire adat_bitclock, // ~12.288 MHz
	input wire oversampling_bitclock, // ~98.304 MHz
	input wire adat_in,
	output wire adat_out,
	output wire[7:0] LED
);

wire data_request;

logic signed [23:0] audio_out [0:7];
adat_out adat_out_0(
        .clk(adat_bitclock),
        .rst(0), .timecode(0), .smux(0),
        .audio_bus(audio_out),
        .adat_bitstream(adat_out),
		  .data_request(data_request)
        );

wire signed [23:0] audio_in [0:7];
wire adat_data_valid;
adat_in adat_in_0(
        .clk(oversampling_bitclock),
        .rst(0),
        .adat_async(adat_in),
        .data_valid(adat_data_valid),
        .audio_bus(audio_in)
        );

logic signed [35:0] dsp_in[8];
wire signed [35:0] dsp_out[8];
int i;
always_comb begin
    for (i=0; i<8; i++) dsp_in[i] <= (audio_in[i] << (36-24));
    for (i=0; i<8; i++) audio_out[i] <= (dsp_out[i] >> (36-24));
end

DSPCore dsp0(
    .clk(oversampling_bitclock),
    .reset(0),
    .start(data_request),
    .inputs(dsp_in),
    .outputs(dsp_out));

wire [23:0] meter_src = audio_out[0];
wire [23:0] abs_val;
assign abs_val = meter_src[23] ? -meter_src : meter_src;

assign LED = abs_val[23:16];

endmodule
